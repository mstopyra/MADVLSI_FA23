magic
tech sky130A
timestamp 1697751355
<< nwell >>
rect -1760 2300 -220 3765
<< nmos >>
rect -1535 920 -1485 2120
rect -1435 920 -1385 2120
rect -1335 920 -1285 2120
rect -1150 920 -1100 2120
rect -880 920 -830 2120
rect -695 920 -645 2120
rect -595 920 -545 2120
rect -495 920 -445 2120
rect -1465 -570 -1415 630
rect -1365 -570 -1315 630
rect -1265 -570 -1215 630
rect -1165 -570 -1115 630
rect -1065 -570 -1015 630
rect -965 -570 -915 630
rect -865 -570 -815 630
rect -765 -570 -715 630
rect -665 -570 -615 630
rect -565 -570 -515 630
<< pmos >>
rect -1465 2410 -1415 3610
rect -1365 2410 -1315 3610
rect -1265 2410 -1215 3610
rect -1165 2410 -1115 3610
rect -1065 2410 -1015 3610
rect -965 2410 -915 3610
rect -865 2410 -815 3610
rect -765 2410 -715 3610
rect -665 2410 -615 3610
rect -565 2410 -515 3610
<< ndiff >>
rect -1585 2105 -1535 2120
rect -1585 935 -1570 2105
rect -1550 935 -1535 2105
rect -1585 920 -1535 935
rect -1485 2105 -1435 2120
rect -1485 935 -1470 2105
rect -1450 935 -1435 2105
rect -1485 920 -1435 935
rect -1385 2105 -1335 2120
rect -1385 935 -1370 2105
rect -1350 935 -1335 2105
rect -1385 920 -1335 935
rect -1285 2105 -1235 2120
rect -1285 935 -1270 2105
rect -1250 935 -1235 2105
rect -1285 920 -1235 935
rect -1200 2105 -1150 2120
rect -1200 935 -1185 2105
rect -1165 935 -1150 2105
rect -1200 920 -1150 935
rect -1100 2105 -1050 2120
rect -1100 935 -1085 2105
rect -1065 935 -1050 2105
rect -1100 920 -1050 935
rect -930 2105 -880 2120
rect -930 935 -915 2105
rect -895 935 -880 2105
rect -930 920 -880 935
rect -830 2105 -780 2120
rect -830 935 -815 2105
rect -795 935 -780 2105
rect -830 920 -780 935
rect -745 2105 -695 2120
rect -745 935 -730 2105
rect -710 935 -695 2105
rect -745 920 -695 935
rect -645 2105 -595 2120
rect -645 935 -630 2105
rect -610 935 -595 2105
rect -645 920 -595 935
rect -545 2105 -495 2120
rect -545 935 -530 2105
rect -510 935 -495 2105
rect -545 920 -495 935
rect -445 2105 -395 2120
rect -445 935 -430 2105
rect -410 935 -395 2105
rect -445 920 -395 935
rect -1515 615 -1465 630
rect -1515 -555 -1500 615
rect -1480 -555 -1465 615
rect -1515 -570 -1465 -555
rect -1415 615 -1365 630
rect -1415 -555 -1400 615
rect -1380 -555 -1365 615
rect -1415 -570 -1365 -555
rect -1315 -570 -1265 630
rect -1215 615 -1165 630
rect -1215 -555 -1200 615
rect -1180 -555 -1165 615
rect -1215 -570 -1165 -555
rect -1115 -570 -1065 630
rect -1015 615 -965 630
rect -1015 -555 -1000 615
rect -980 -555 -965 615
rect -1015 -570 -965 -555
rect -915 -570 -865 630
rect -815 615 -765 630
rect -815 -555 -800 615
rect -780 -555 -765 615
rect -815 -570 -765 -555
rect -715 -570 -665 630
rect -615 615 -565 630
rect -615 -555 -600 615
rect -580 -555 -565 615
rect -615 -570 -565 -555
rect -515 615 -465 630
rect -515 -555 -500 615
rect -480 -555 -465 615
rect -515 -570 -465 -555
<< pdiff >>
rect -1515 3595 -1465 3610
rect -1515 2425 -1500 3595
rect -1480 2425 -1465 3595
rect -1515 2410 -1465 2425
rect -1415 3595 -1365 3610
rect -1415 2425 -1400 3595
rect -1380 2425 -1365 3595
rect -1415 2410 -1365 2425
rect -1315 3595 -1265 3610
rect -1315 2425 -1300 3595
rect -1280 2425 -1265 3595
rect -1315 2410 -1265 2425
rect -1215 3595 -1165 3610
rect -1215 2425 -1200 3595
rect -1180 2425 -1165 3595
rect -1215 2410 -1165 2425
rect -1115 3595 -1065 3610
rect -1115 2425 -1100 3595
rect -1080 2425 -1065 3595
rect -1115 2410 -1065 2425
rect -1015 3595 -965 3610
rect -1015 2425 -1000 3595
rect -980 2425 -965 3595
rect -1015 2410 -965 2425
rect -915 3595 -865 3610
rect -915 2425 -900 3595
rect -880 2425 -865 3595
rect -915 2410 -865 2425
rect -815 3595 -765 3610
rect -815 2425 -800 3595
rect -780 2425 -765 3595
rect -815 2410 -765 2425
rect -715 3595 -665 3610
rect -715 2425 -700 3595
rect -680 2425 -665 3595
rect -715 2410 -665 2425
rect -615 3595 -565 3610
rect -615 2425 -600 3595
rect -580 2425 -565 3595
rect -615 2410 -565 2425
rect -515 3595 -465 3610
rect -515 2425 -500 3595
rect -480 2425 -465 3595
rect -515 2410 -465 2425
<< ndiffc >>
rect -1570 935 -1550 2105
rect -1470 935 -1450 2105
rect -1370 935 -1350 2105
rect -1270 935 -1250 2105
rect -1185 935 -1165 2105
rect -1085 935 -1065 2105
rect -915 935 -895 2105
rect -815 935 -795 2105
rect -730 935 -710 2105
rect -630 935 -610 2105
rect -530 935 -510 2105
rect -430 935 -410 2105
rect -1500 -555 -1480 615
rect -1400 -555 -1380 615
rect -1200 -555 -1180 615
rect -1000 -555 -980 615
rect -800 -555 -780 615
rect -600 -555 -580 615
rect -500 -555 -480 615
<< pdiffc >>
rect -1500 2425 -1480 3595
rect -1400 2425 -1380 3595
rect -1300 2425 -1280 3595
rect -1200 2425 -1180 3595
rect -1100 2425 -1080 3595
rect -1000 2425 -980 3595
rect -900 2425 -880 3595
rect -800 2425 -780 3595
rect -700 2425 -680 3595
rect -600 2425 -580 3595
rect -500 2425 -480 3595
<< psubdiff >>
rect -1635 2105 -1585 2120
rect -1635 935 -1615 2105
rect -1595 935 -1585 2105
rect -1635 920 -1585 935
rect -395 2105 -345 2120
rect -395 935 -380 2105
rect -360 935 -345 2105
rect -395 920 -345 935
rect -465 615 -415 630
rect -465 -555 -450 615
rect -430 -555 -415 615
rect -465 -570 -415 -555
<< nsubdiff >>
rect -1565 3595 -1515 3610
rect -1565 2425 -1550 3595
rect -1530 2425 -1515 3595
rect -1565 2410 -1515 2425
rect -465 3595 -415 3610
rect -465 2425 -450 3595
rect -430 2425 -415 3595
rect -465 2410 -415 2425
<< psubdiffcont >>
rect -1615 935 -1595 2105
rect -380 935 -360 2105
rect -450 -555 -430 615
<< nsubdiffcont >>
rect -1550 2425 -1530 3595
rect -450 2425 -430 3595
<< poly >>
rect -765 3755 -715 3765
rect -765 3725 -755 3755
rect -725 3725 -715 3755
rect -765 3715 -715 3725
rect -1465 3665 -1415 3675
rect -1465 3635 -1455 3665
rect -1425 3635 -1415 3665
rect -1465 3610 -1415 3635
rect -1265 3665 -715 3715
rect -1365 3610 -1315 3625
rect -1265 3610 -1215 3665
rect -1165 3610 -1115 3665
rect -1065 3610 -1015 3625
rect -965 3610 -915 3625
rect -865 3610 -815 3665
rect -765 3610 -715 3665
rect -565 3665 -515 3675
rect -565 3635 -555 3665
rect -525 3635 -515 3665
rect -665 3610 -615 3625
rect -565 3610 -515 3635
rect -1465 2395 -1415 2410
rect -1365 2370 -1315 2410
rect -1265 2395 -1215 2410
rect -1165 2395 -1115 2410
rect -1065 2370 -1015 2410
rect -965 2370 -915 2410
rect -865 2395 -815 2410
rect -765 2395 -715 2410
rect -665 2370 -615 2410
rect -565 2395 -515 2410
rect -1365 2360 -220 2370
rect -1365 2330 -260 2360
rect -230 2330 -220 2360
rect -1365 2320 -220 2330
rect -1760 2270 -1095 2280
rect -1760 2240 -1750 2270
rect -1720 2240 -1095 2270
rect -1760 2230 -1095 2240
rect -1155 2225 -1095 2230
rect -1150 2185 -1095 2225
rect -695 2275 -220 2285
rect -695 2245 -260 2275
rect -230 2245 -220 2275
rect -695 2235 -220 2245
rect -1150 2135 -830 2185
rect -1535 2120 -1485 2135
rect -1435 2120 -1385 2135
rect -1335 2120 -1285 2135
rect -1150 2120 -1100 2135
rect -880 2120 -830 2135
rect -695 2120 -645 2235
rect -595 2120 -545 2135
rect -495 2120 -445 2135
rect -1535 895 -1485 920
rect -1535 865 -1525 895
rect -1495 865 -1485 895
rect -1535 855 -1485 865
rect -1435 800 -1385 920
rect -1335 880 -1285 920
rect -1150 905 -1100 920
rect -880 905 -830 920
rect -695 880 -645 920
rect -1335 830 -645 880
rect -595 800 -545 920
rect -495 895 -445 920
rect -495 865 -485 895
rect -455 865 -445 895
rect -495 855 -445 865
rect -1760 790 -545 800
rect -1760 760 -1750 790
rect -1720 760 -545 790
rect -1760 750 -545 760
rect -1365 710 -220 720
rect -1365 680 -260 710
rect -230 680 -220 710
rect -1365 670 -220 680
rect -1465 630 -1415 645
rect -1365 630 -1315 670
rect -1265 630 -1215 645
rect -1165 630 -1115 645
rect -1065 630 -1015 670
rect -965 630 -915 670
rect -865 630 -815 645
rect -765 630 -715 645
rect -665 630 -615 670
rect -565 630 -515 645
rect -1465 -635 -1415 -570
rect -1365 -585 -1315 -570
rect -1265 -585 -1215 -570
rect -1165 -585 -1115 -570
rect -1065 -585 -1015 -570
rect -965 -585 -915 -570
rect -865 -585 -815 -570
rect -765 -585 -715 -570
rect -665 -585 -615 -570
rect -1265 -595 -1115 -585
rect -1265 -625 -1255 -595
rect -1225 -625 -1115 -595
rect -1265 -635 -1115 -625
rect -865 -595 -715 -585
rect -865 -625 -755 -595
rect -725 -625 -715 -595
rect -865 -635 -715 -625
rect -1520 -645 -1415 -635
rect -1520 -675 -1510 -645
rect -1480 -675 -1415 -645
rect -1520 -685 -1415 -675
rect -565 -645 -515 -570
rect -565 -655 -460 -645
rect -565 -685 -500 -655
rect -470 -685 -460 -655
rect -565 -695 -460 -685
<< polycont >>
rect -755 3725 -725 3755
rect -1455 3635 -1425 3665
rect -555 3635 -525 3665
rect -260 2330 -230 2360
rect -1750 2240 -1720 2270
rect -260 2245 -230 2275
rect -1525 865 -1495 895
rect -485 865 -455 895
rect -1750 760 -1720 790
rect -260 680 -230 710
rect -1255 -625 -1225 -595
rect -755 -625 -725 -595
rect -1510 -675 -1480 -645
rect -500 -685 -470 -655
<< locali >>
rect -890 3755 -715 3765
rect -890 3725 -755 3755
rect -725 3725 -715 3755
rect -890 3715 -715 3725
rect -1515 3665 -1415 3675
rect -1515 3635 -1455 3665
rect -1425 3635 -1415 3665
rect -1515 3625 -1415 3635
rect -565 3665 -470 3675
rect -565 3635 -555 3665
rect -525 3635 -470 3665
rect -565 3625 -470 3635
rect -1515 3605 -1470 3625
rect -510 3605 -470 3625
rect -1560 3595 -1470 3605
rect -1560 2425 -1550 3595
rect -1530 2425 -1500 3595
rect -1480 2425 -1470 3595
rect -1560 2415 -1470 2425
rect -1410 3595 -1370 3605
rect -1410 2425 -1400 3595
rect -1380 2425 -1370 3595
rect -1410 2385 -1370 2425
rect -1690 2345 -1370 2385
rect -1310 3595 -1270 3605
rect -1310 2425 -1300 3595
rect -1280 2425 -1270 3595
rect -1760 2270 -1710 2280
rect -1760 2240 -1750 2270
rect -1720 2240 -1710 2270
rect -1760 2115 -1710 2240
rect -1760 790 -1710 915
rect -1760 760 -1750 790
rect -1720 760 -1710 790
rect -1760 750 -1710 760
rect -1690 725 -1650 2345
rect -1310 2285 -1270 2425
rect -1210 3595 -1170 3605
rect -1210 2425 -1200 3595
rect -1180 2425 -1170 3595
rect -1210 2415 -1170 2425
rect -1110 3595 -1070 3605
rect -1110 2425 -1100 3595
rect -1080 2425 -1070 3595
rect -1480 2245 -1270 2285
rect -1110 2285 -1070 2425
rect -1010 3595 -970 3605
rect -1010 2425 -1000 3595
rect -980 2425 -970 3595
rect -1110 2255 -1055 2285
rect -1630 2105 -1540 2115
rect -1630 935 -1615 2105
rect -1595 935 -1570 2105
rect -1550 935 -1540 2105
rect -1630 925 -1540 935
rect -1480 2105 -1440 2245
rect -1480 935 -1470 2105
rect -1450 935 -1440 2105
rect -1480 925 -1440 935
rect -1380 2160 -1155 2200
rect -1380 2105 -1340 2160
rect -1380 935 -1370 2105
rect -1350 935 -1340 2105
rect -1380 925 -1340 935
rect -1280 2105 -1240 2115
rect -1280 935 -1270 2105
rect -1250 935 -1240 2105
rect -1585 905 -1540 925
rect -1585 895 -1485 905
rect -1585 865 -1525 895
rect -1495 865 -1485 895
rect -1585 855 -1485 865
rect -1690 685 -1370 725
rect -1510 615 -1470 625
rect -1510 -555 -1500 615
rect -1480 -555 -1470 615
rect -1510 -635 -1470 -555
rect -1410 615 -1370 685
rect -1280 720 -1240 935
rect -1195 2105 -1155 2160
rect -1195 935 -1185 2105
rect -1165 935 -1155 2105
rect -1195 925 -1155 935
rect -1095 2105 -1055 2255
rect -1095 935 -1085 2105
rect -1065 935 -1055 2105
rect -1095 925 -1055 935
rect -1280 680 -1170 720
rect -1410 -555 -1400 615
rect -1380 -555 -1370 615
rect -1410 -595 -1370 -555
rect -1210 615 -1170 680
rect -1210 -555 -1200 615
rect -1180 -555 -1170 615
rect -1210 -565 -1170 -555
rect -1010 615 -970 2425
rect -910 3595 -870 3605
rect -910 2425 -900 3595
rect -880 2425 -870 3595
rect -910 2285 -870 2425
rect -810 3595 -770 3605
rect -810 2425 -800 3595
rect -780 2425 -770 3595
rect -810 2415 -770 2425
rect -710 3595 -670 3605
rect -710 2425 -700 3595
rect -680 2425 -670 3595
rect -925 2245 -870 2285
rect -710 2275 -670 2425
rect -610 3595 -570 3605
rect -610 2425 -600 3595
rect -580 2425 -570 3595
rect -610 2380 -570 2425
rect -510 3595 -420 3605
rect -510 2425 -500 3595
rect -480 2425 -450 3595
rect -430 2425 -420 3595
rect -510 2415 -420 2425
rect -610 2340 -290 2380
rect -925 2105 -885 2245
rect -710 2235 -500 2275
rect -925 935 -915 2105
rect -895 935 -885 2105
rect -925 925 -885 935
rect -825 2160 -600 2200
rect -825 2105 -785 2160
rect -825 935 -815 2105
rect -795 935 -785 2105
rect -825 925 -785 935
rect -740 2105 -700 2115
rect -740 935 -730 2105
rect -710 935 -700 2105
rect -740 720 -700 935
rect -640 2105 -600 2160
rect -640 935 -630 2105
rect -610 935 -600 2105
rect -640 925 -600 935
rect -540 2105 -500 2235
rect -540 935 -530 2105
rect -510 935 -500 2105
rect -540 925 -500 935
rect -440 2105 -350 2115
rect -440 935 -430 2105
rect -410 935 -380 2105
rect -360 935 -350 2105
rect -440 925 -350 935
rect -440 905 -395 925
rect -495 895 -395 905
rect -495 865 -485 895
rect -455 865 -395 895
rect -495 855 -395 865
rect -330 790 -290 2340
rect -270 2360 -220 2485
rect -270 2330 -260 2360
rect -230 2330 -220 2360
rect -270 2320 -220 2330
rect -270 2275 -220 2285
rect -270 2245 -260 2275
rect -230 2245 -220 2275
rect -270 2120 -220 2245
rect -1010 -555 -1000 615
rect -980 -555 -970 615
rect -1265 -595 -1215 -585
rect -1410 -625 -1255 -595
rect -1225 -625 -1215 -595
rect -1410 -635 -1215 -625
rect -1520 -645 -1470 -635
rect -1520 -675 -1510 -645
rect -1480 -675 -1470 -645
rect -1520 -685 -1470 -675
rect -1010 -680 -970 -555
rect -810 680 -700 720
rect -610 750 -290 790
rect -810 615 -770 680
rect -810 -555 -800 615
rect -780 -555 -770 615
rect -810 -565 -770 -555
rect -610 615 -570 750
rect -270 710 -220 720
rect -270 680 -260 710
rect -230 680 -220 710
rect -610 -555 -600 615
rect -580 -555 -570 615
rect -765 -595 -715 -585
rect -610 -595 -570 -555
rect -765 -625 -755 -595
rect -725 -625 -570 -595
rect -765 -635 -570 -625
rect -510 615 -420 625
rect -510 -555 -500 615
rect -480 -555 -450 615
rect -430 -555 -420 615
rect -270 555 -220 680
rect -510 -565 -420 -555
rect -510 -645 -470 -565
rect -510 -655 -460 -645
rect -1050 -730 -935 -680
rect -510 -685 -500 -655
rect -470 -685 -460 -655
rect -510 -695 -460 -685
<< viali >>
rect -1550 2800 -1530 3375
rect -1500 2800 -1480 3375
rect -1200 2800 -1180 3375
rect -1615 1195 -1595 1770
rect -1570 1195 -1550 1770
rect -1270 1195 -1250 1770
rect -1500 -270 -1480 305
rect -1200 -265 -1180 310
rect -800 2805 -780 3380
rect -500 2800 -480 3375
rect -450 2800 -430 3375
rect -730 1195 -710 1770
rect -430 1200 -410 1775
rect -380 1195 -360 1770
rect -800 -265 -780 310
rect -500 -260 -480 315
rect -450 -265 -430 310
<< metal1 >>
rect -1760 3380 -220 3385
rect -1760 3375 -800 3380
rect -1760 2800 -1550 3375
rect -1530 2800 -1500 3375
rect -1480 2800 -1200 3375
rect -1180 2805 -800 3375
rect -780 3375 -220 3380
rect -780 2805 -500 3375
rect -1180 2800 -500 2805
rect -480 2800 -450 3375
rect -430 2800 -220 3375
rect -1760 2790 -220 2800
rect -1760 1775 -220 1780
rect -1760 1770 -430 1775
rect -1760 1195 -1615 1770
rect -1595 1195 -1570 1770
rect -1550 1195 -1270 1770
rect -1250 1195 -730 1770
rect -710 1200 -430 1770
rect -410 1770 -220 1775
rect -410 1200 -380 1770
rect -710 1195 -380 1200
rect -360 1195 -220 1770
rect -1760 1185 -220 1195
rect -1760 315 -220 320
rect -1760 310 -500 315
rect -1760 305 -1200 310
rect -1760 -270 -1500 305
rect -1480 -265 -1200 305
rect -1180 -265 -800 310
rect -780 -260 -500 310
rect -480 310 -220 315
rect -480 -260 -450 310
rect -780 -265 -450 -260
rect -430 -265 -220 310
rect -1480 -270 -220 -265
rect -1760 -275 -220 -270
<< labels >>
rlabel locali -810 3765 -810 3765 1 VBP
rlabel metal1 -1760 3075 -1760 3075 7 VDD
rlabel locali -1760 2185 -1760 2185 7 V2
rlabel metal1 -1760 1480 -1760 1480 7 GND
rlabel locali -1760 845 -1760 845 7 V1
rlabel metal1 -1760 -5 -1760 -5 7 GND
rlabel locali -990 -730 -990 -730 5 VOUT
rlabel locali -220 625 -220 625 3 VCN
rlabel locali -220 2185 -220 2185 3 VBN
rlabel locali -220 2415 -220 2415 3 VCP
<< end >>
