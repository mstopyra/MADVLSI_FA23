magic
tech sky130A
timestamp 1697397656
<< nwell >>
rect -2415 -145 -930 1300
rect -2435 -4035 -1115 -2250
<< nmos >>
rect -2330 -1470 -2280 -270
rect -2225 -1470 -2175 -270
rect -2150 -1470 -2100 -270
rect -2075 -1470 -2025 -270
rect -2000 -1470 -1950 -270
rect -1925 -1470 -1875 -270
rect -1820 -1470 -1770 -270
rect -1745 -1470 -1695 -270
rect -1670 -1470 -1620 -270
rect -1595 -1470 -1545 -270
rect -1520 -1470 -1470 -270
rect -1305 -1470 -1255 -270
rect -2370 -1735 -1170 -1685
rect -2370 -1950 -1170 -1900
rect -2370 -2055 -1170 -2005
rect -2370 -2160 -1170 -2110
rect -2335 -5375 -2285 -4175
rect -2230 -5375 -2180 -4175
rect -2125 -5375 -2075 -4175
rect -2020 -5375 -1970 -4175
rect -1915 -5375 -1865 -4175
rect -1810 -5375 -1760 -4175
rect -1595 -5375 -1545 -4175
rect -1490 -5375 -1440 -4175
rect -1385 -5375 -1335 -4175
rect -1280 -5375 -1230 -4175
rect -1175 -5375 -1125 -4175
rect -1070 -5375 -1020 -4175
<< pmos >>
rect -2330 -90 -2280 1110
rect -2225 -90 -2175 1110
rect -2120 -90 -2070 1110
rect -2015 -90 -1965 1110
rect -1910 -90 -1860 1110
rect -1805 -90 -1755 1110
rect -1590 -90 -1540 1110
rect -1485 -90 -1435 1110
rect -1380 -90 -1330 1110
rect -1275 -90 -1225 1110
rect -1170 -90 -1120 1110
rect -1065 -90 -1015 1110
rect -2370 -2375 -1170 -2325
rect -2370 -2590 -1170 -2540
rect -2335 -3995 -2285 -2795
rect -2230 -3995 -2180 -2795
rect -2155 -3995 -2105 -2795
rect -2080 -3995 -2030 -2795
rect -2005 -3995 -1955 -2795
rect -1930 -3995 -1880 -2795
rect -1825 -3995 -1775 -2795
rect -1750 -3995 -1700 -2795
rect -1675 -3995 -1625 -2795
rect -1600 -3995 -1550 -2795
rect -1525 -3995 -1475 -2795
rect -1310 -3995 -1260 -2795
<< ndiff >>
rect -2385 -285 -2330 -270
rect -2385 -1455 -2370 -285
rect -2345 -1455 -2330 -285
rect -2385 -1470 -2330 -1455
rect -2280 -285 -2225 -270
rect -2280 -1455 -2265 -285
rect -2240 -1455 -2225 -285
rect -2280 -1470 -2225 -1455
rect -2175 -1470 -2150 -270
rect -2100 -1470 -2075 -270
rect -2025 -1470 -2000 -270
rect -1950 -1470 -1925 -270
rect -1875 -285 -1820 -270
rect -1875 -1455 -1860 -285
rect -1835 -1455 -1820 -285
rect -1875 -1470 -1820 -1455
rect -1770 -1470 -1745 -270
rect -1695 -1470 -1670 -270
rect -1620 -1470 -1595 -270
rect -1545 -1470 -1520 -270
rect -1470 -285 -1415 -270
rect -1360 -285 -1305 -270
rect -1470 -1455 -1455 -285
rect -1430 -1455 -1415 -285
rect -1360 -1455 -1345 -285
rect -1320 -1455 -1305 -285
rect -1470 -1470 -1415 -1455
rect -1360 -1470 -1305 -1455
rect -1255 -285 -1200 -270
rect -1255 -1455 -1240 -285
rect -1215 -1455 -1200 -285
rect -1255 -1470 -1200 -1455
rect -2370 -1645 -1170 -1630
rect -2370 -1670 -2355 -1645
rect -1185 -1670 -1170 -1645
rect -2370 -1685 -1170 -1670
rect -2370 -1750 -1170 -1735
rect -2370 -1775 -2355 -1750
rect -1185 -1775 -1170 -1750
rect -2370 -1790 -1170 -1775
rect -2370 -1860 -1170 -1845
rect -2370 -1885 -2355 -1860
rect -1185 -1885 -1170 -1860
rect -2370 -1900 -1170 -1885
rect -2370 -1965 -1170 -1950
rect -2370 -1990 -2355 -1965
rect -1185 -1990 -1170 -1965
rect -2370 -2005 -1170 -1990
rect -2370 -2070 -1170 -2055
rect -2370 -2095 -2355 -2070
rect -1185 -2095 -1170 -2070
rect -2370 -2110 -1170 -2095
rect -2370 -2175 -1170 -2160
rect -2370 -2200 -2355 -2175
rect -1185 -2200 -1170 -2175
rect -2370 -2215 -1170 -2200
rect -2390 -4190 -2335 -4175
rect -2390 -5360 -2375 -4190
rect -2350 -5360 -2335 -4190
rect -2390 -5375 -2335 -5360
rect -2285 -4190 -2230 -4175
rect -2285 -5360 -2270 -4190
rect -2245 -5360 -2230 -4190
rect -2285 -5375 -2230 -5360
rect -2180 -4190 -2125 -4175
rect -2180 -5360 -2165 -4190
rect -2140 -5360 -2125 -4190
rect -2180 -5375 -2125 -5360
rect -2075 -4190 -2020 -4175
rect -2075 -5360 -2060 -4190
rect -2035 -5360 -2020 -4190
rect -2075 -5375 -2020 -5360
rect -1970 -4190 -1915 -4175
rect -1970 -5360 -1955 -4190
rect -1930 -5360 -1915 -4190
rect -1970 -5375 -1915 -5360
rect -1865 -4190 -1810 -4175
rect -1865 -5360 -1850 -4190
rect -1825 -5360 -1810 -4190
rect -1865 -5375 -1810 -5360
rect -1760 -4190 -1705 -4175
rect -1650 -4190 -1595 -4175
rect -1760 -5360 -1745 -4190
rect -1720 -5360 -1705 -4190
rect -1650 -5360 -1635 -4190
rect -1610 -5360 -1595 -4190
rect -1760 -5375 -1705 -5360
rect -1650 -5375 -1595 -5360
rect -1545 -4190 -1490 -4175
rect -1545 -5360 -1530 -4190
rect -1505 -5360 -1490 -4190
rect -1545 -5375 -1490 -5360
rect -1440 -4190 -1385 -4175
rect -1440 -5360 -1425 -4190
rect -1400 -5360 -1385 -4190
rect -1440 -5375 -1385 -5360
rect -1335 -4190 -1280 -4175
rect -1335 -5360 -1320 -4190
rect -1295 -5360 -1280 -4190
rect -1335 -5375 -1280 -5360
rect -1230 -4190 -1175 -4175
rect -1230 -5360 -1215 -4190
rect -1190 -5360 -1175 -4190
rect -1230 -5375 -1175 -5360
rect -1125 -4190 -1070 -4175
rect -1125 -5360 -1110 -4190
rect -1085 -5360 -1070 -4190
rect -1125 -5375 -1070 -5360
rect -1020 -4190 -965 -4175
rect -1020 -5360 -1005 -4190
rect -980 -5360 -965 -4190
rect -1020 -5375 -965 -5360
<< pdiff >>
rect -2385 1095 -2330 1110
rect -2385 -75 -2370 1095
rect -2345 -75 -2330 1095
rect -2385 -90 -2330 -75
rect -2280 1095 -2225 1110
rect -2280 -75 -2265 1095
rect -2240 -75 -2225 1095
rect -2280 -90 -2225 -75
rect -2175 1095 -2120 1110
rect -2175 -75 -2160 1095
rect -2135 -75 -2120 1095
rect -2175 -90 -2120 -75
rect -2070 1095 -2015 1110
rect -2070 -75 -2055 1095
rect -2030 -75 -2015 1095
rect -2070 -90 -2015 -75
rect -1965 1095 -1910 1110
rect -1965 -75 -1950 1095
rect -1925 -75 -1910 1095
rect -1965 -90 -1910 -75
rect -1860 1095 -1805 1110
rect -1860 -75 -1845 1095
rect -1820 -75 -1805 1095
rect -1860 -90 -1805 -75
rect -1755 1095 -1700 1110
rect -1645 1095 -1590 1110
rect -1755 -75 -1740 1095
rect -1715 -75 -1700 1095
rect -1645 -75 -1630 1095
rect -1605 -75 -1590 1095
rect -1755 -90 -1700 -75
rect -1645 -90 -1590 -75
rect -1540 1095 -1485 1110
rect -1540 -75 -1525 1095
rect -1500 -75 -1485 1095
rect -1540 -90 -1485 -75
rect -1435 1095 -1380 1110
rect -1435 -75 -1420 1095
rect -1395 -75 -1380 1095
rect -1435 -90 -1380 -75
rect -1330 1095 -1275 1110
rect -1330 -75 -1315 1095
rect -1290 -75 -1275 1095
rect -1330 -90 -1275 -75
rect -1225 1095 -1170 1110
rect -1225 -75 -1210 1095
rect -1185 -75 -1170 1095
rect -1225 -90 -1170 -75
rect -1120 1095 -1065 1110
rect -1120 -75 -1105 1095
rect -1080 -75 -1065 1095
rect -1120 -90 -1065 -75
rect -1015 1095 -960 1110
rect -1015 -75 -1000 1095
rect -975 -75 -960 1095
rect -1015 -90 -960 -75
rect -2370 -2285 -1170 -2270
rect -2370 -2310 -2355 -2285
rect -1185 -2310 -1170 -2285
rect -2370 -2325 -1170 -2310
rect -2370 -2390 -1170 -2375
rect -2370 -2415 -2355 -2390
rect -1185 -2415 -1170 -2390
rect -2370 -2430 -1170 -2415
rect -2370 -2500 -1170 -2485
rect -2370 -2525 -2355 -2500
rect -1185 -2525 -1170 -2500
rect -2370 -2540 -1170 -2525
rect -2370 -2605 -1170 -2590
rect -2370 -2630 -2355 -2605
rect -1185 -2630 -1170 -2605
rect -2370 -2645 -1170 -2630
rect -2390 -2810 -2335 -2795
rect -2390 -3980 -2375 -2810
rect -2350 -3980 -2335 -2810
rect -2390 -3995 -2335 -3980
rect -2285 -2810 -2230 -2795
rect -2285 -3980 -2270 -2810
rect -2245 -3980 -2230 -2810
rect -2285 -3995 -2230 -3980
rect -2180 -3995 -2155 -2795
rect -2105 -3995 -2080 -2795
rect -2030 -3995 -2005 -2795
rect -1955 -3995 -1930 -2795
rect -1880 -2810 -1825 -2795
rect -1880 -3980 -1865 -2810
rect -1840 -3980 -1825 -2810
rect -1880 -3995 -1825 -3980
rect -1775 -3995 -1750 -2795
rect -1700 -3995 -1675 -2795
rect -1625 -3995 -1600 -2795
rect -1550 -3995 -1525 -2795
rect -1475 -2810 -1420 -2795
rect -1365 -2810 -1310 -2795
rect -1475 -3980 -1460 -2810
rect -1435 -3980 -1420 -2810
rect -1365 -3980 -1350 -2810
rect -1325 -3980 -1310 -2810
rect -1475 -3995 -1420 -3980
rect -1365 -3995 -1310 -3980
rect -1260 -2810 -1205 -2795
rect -1260 -3980 -1245 -2810
rect -1220 -3980 -1205 -2810
rect -1260 -3995 -1205 -3980
<< ndiffc >>
rect -2370 -1455 -2345 -285
rect -2265 -1455 -2240 -285
rect -1860 -1455 -1835 -285
rect -1455 -1455 -1430 -285
rect -1345 -1455 -1320 -285
rect -1240 -1455 -1215 -285
rect -2355 -1670 -1185 -1645
rect -2355 -1775 -1185 -1750
rect -2355 -1885 -1185 -1860
rect -2355 -1990 -1185 -1965
rect -2355 -2095 -1185 -2070
rect -2355 -2200 -1185 -2175
rect -2375 -5360 -2350 -4190
rect -2270 -5360 -2245 -4190
rect -2165 -5360 -2140 -4190
rect -2060 -5360 -2035 -4190
rect -1955 -5360 -1930 -4190
rect -1850 -5360 -1825 -4190
rect -1745 -5360 -1720 -4190
rect -1635 -5360 -1610 -4190
rect -1530 -5360 -1505 -4190
rect -1425 -5360 -1400 -4190
rect -1320 -5360 -1295 -4190
rect -1215 -5360 -1190 -4190
rect -1110 -5360 -1085 -4190
rect -1005 -5360 -980 -4190
<< pdiffc >>
rect -2370 -75 -2345 1095
rect -2265 -75 -2240 1095
rect -2160 -75 -2135 1095
rect -2055 -75 -2030 1095
rect -1950 -75 -1925 1095
rect -1845 -75 -1820 1095
rect -1740 -75 -1715 1095
rect -1630 -75 -1605 1095
rect -1525 -75 -1500 1095
rect -1420 -75 -1395 1095
rect -1315 -75 -1290 1095
rect -1210 -75 -1185 1095
rect -1105 -75 -1080 1095
rect -1000 -75 -975 1095
rect -2355 -2310 -1185 -2285
rect -2355 -2415 -1185 -2390
rect -2355 -2525 -1185 -2500
rect -2355 -2630 -1185 -2605
rect -2375 -3980 -2350 -2810
rect -2270 -3980 -2245 -2810
rect -1865 -3980 -1840 -2810
rect -1460 -3980 -1435 -2810
rect -1350 -3980 -1325 -2810
rect -1245 -3980 -1220 -2810
<< psubdiff >>
rect -1415 -285 -1360 -270
rect -1415 -1455 -1400 -285
rect -1375 -1455 -1360 -285
rect -1415 -1470 -1360 -1455
rect -2370 -1805 -1170 -1790
rect -2370 -1830 -2355 -1805
rect -1185 -1830 -1170 -1805
rect -2370 -1845 -1170 -1830
rect -1705 -4190 -1650 -4175
rect -1705 -5360 -1690 -4190
rect -1665 -5360 -1650 -4190
rect -1705 -5375 -1650 -5360
<< nsubdiff >>
rect -1700 1095 -1645 1110
rect -1700 -75 -1685 1095
rect -1660 -75 -1645 1095
rect -1700 -90 -1645 -75
rect -2370 -2445 -1170 -2430
rect -2370 -2470 -2355 -2445
rect -1185 -2470 -1170 -2445
rect -2370 -2485 -1170 -2470
rect -1420 -2810 -1365 -2795
rect -1420 -3980 -1405 -2810
rect -1380 -3980 -1365 -2810
rect -1420 -3995 -1365 -3980
<< psubdiffcont >>
rect -1400 -1455 -1375 -285
rect -2355 -1830 -1185 -1805
rect -1690 -5360 -1665 -4190
<< nsubdiffcont >>
rect -1685 -75 -1660 1095
rect -2355 -2470 -1185 -2445
rect -1405 -3980 -1380 -2810
<< poly >>
rect -2330 1110 -2280 1125
rect -2225 1110 -2175 1125
rect -2120 1110 -2070 1125
rect -2015 1110 -1965 1125
rect -1910 1110 -1860 1125
rect -1805 1110 -1755 1125
rect -1590 1110 -1540 1125
rect -1485 1110 -1435 1125
rect -1380 1110 -1330 1125
rect -1275 1110 -1225 1125
rect -1170 1110 -1120 1125
rect -1065 1110 -1015 1125
rect -2330 -160 -2280 -90
rect -2225 -105 -2175 -90
rect -2120 -105 -2070 -90
rect -2015 -105 -1965 -90
rect -1910 -105 -1860 -90
rect -1805 -105 -1755 -90
rect -1590 -105 -1540 -90
rect -1485 -105 -1435 -90
rect -1380 -105 -1330 -90
rect -1275 -105 -1225 -90
rect -1170 -105 -1120 -90
rect -2225 -115 -1120 -105
rect -2225 -145 -2165 -115
rect -2130 -145 -2060 -115
rect -2025 -145 -1955 -115
rect -1920 -145 -1745 -115
rect -1710 -145 -1425 -115
rect -1390 -145 -1320 -115
rect -1285 -145 -1215 -115
rect -1180 -145 -1120 -115
rect -2225 -155 -1120 -145
rect -2380 -170 -2280 -160
rect -2380 -200 -2370 -170
rect -2340 -200 -2280 -170
rect -1065 -180 -1015 -90
rect -2380 -210 -2280 -200
rect -1125 -190 -1015 -180
rect -1125 -220 -1115 -190
rect -1085 -220 -1015 -190
rect -1125 -230 -1015 -220
rect -2330 -270 -2280 -255
rect -2225 -270 -2175 -255
rect -2150 -270 -2100 -255
rect -2075 -270 -2025 -255
rect -2000 -270 -1950 -255
rect -1925 -270 -1875 -255
rect -1820 -270 -1770 -255
rect -1745 -270 -1695 -255
rect -1670 -270 -1620 -255
rect -1595 -270 -1545 -255
rect -1520 -270 -1470 -255
rect -1305 -270 -1255 -255
rect -2330 -1485 -2280 -1470
rect -2225 -1485 -2175 -1470
rect -2150 -1485 -2100 -1470
rect -2075 -1485 -2025 -1470
rect -2000 -1485 -1950 -1470
rect -1925 -1485 -1875 -1470
rect -1820 -1485 -1770 -1470
rect -1745 -1485 -1695 -1470
rect -1670 -1485 -1620 -1470
rect -1595 -1485 -1545 -1470
rect -1520 -1485 -1470 -1470
rect -1305 -1485 -1255 -1470
rect -2440 -1535 -1255 -1485
rect -2440 -1645 -2390 -1535
rect -2440 -1675 -2430 -1645
rect -2400 -1675 -2390 -1645
rect -2440 -1685 -2390 -1675
rect -2440 -1735 -2370 -1685
rect -1170 -1735 -1155 -1685
rect -2440 -1900 -2385 -1735
rect -2440 -1950 -2370 -1900
rect -1170 -1950 -1155 -1900
rect -2440 -2005 -2385 -1950
rect -2440 -2055 -2370 -2005
rect -1170 -2055 -1155 -2005
rect -2440 -2110 -2385 -2055
rect -2440 -2160 -2370 -2110
rect -1170 -2120 -1105 -2110
rect -1170 -2150 -1145 -2120
rect -1115 -2150 -1105 -2120
rect -1170 -2160 -1105 -2150
rect -2385 -2375 -2370 -2325
rect -1170 -2375 -1155 -2325
rect -2385 -2590 -2370 -2540
rect -1170 -2590 -1155 -2540
rect -2335 -2690 -2285 -2680
rect -2335 -2720 -2325 -2690
rect -2295 -2720 -2285 -2690
rect -2335 -2730 -2285 -2720
rect -2335 -2780 -1260 -2730
rect -2335 -2795 -2285 -2780
rect -2230 -2795 -2180 -2780
rect -2155 -2795 -2105 -2780
rect -2080 -2795 -2030 -2780
rect -2005 -2795 -1955 -2780
rect -1930 -2795 -1880 -2780
rect -1825 -2795 -1775 -2780
rect -1750 -2795 -1700 -2780
rect -1675 -2795 -1625 -2780
rect -1600 -2795 -1550 -2780
rect -1525 -2795 -1475 -2780
rect -1310 -2795 -1260 -2780
rect -2335 -4010 -2285 -3995
rect -2230 -4010 -2180 -3995
rect -2155 -4010 -2105 -3995
rect -2080 -4010 -2030 -3995
rect -2005 -4010 -1955 -3995
rect -1930 -4010 -1880 -3995
rect -1825 -4010 -1775 -3995
rect -1750 -4010 -1700 -3995
rect -1675 -4010 -1625 -3995
rect -1600 -4010 -1550 -3995
rect -1525 -4010 -1475 -3995
rect -1310 -4010 -1260 -3995
rect -1130 -4045 -1020 -4035
rect -2385 -4065 -2285 -4055
rect -2385 -4095 -2375 -4065
rect -2345 -4095 -2285 -4065
rect -1130 -4075 -1120 -4045
rect -1090 -4075 -1020 -4045
rect -1130 -4085 -1020 -4075
rect -2385 -4105 -2285 -4095
rect -2335 -4175 -2285 -4105
rect -2230 -4120 -1125 -4110
rect -2230 -4150 -2170 -4120
rect -2135 -4150 -2065 -4120
rect -2030 -4150 -1960 -4120
rect -1925 -4150 -1750 -4120
rect -1715 -4150 -1430 -4120
rect -1395 -4150 -1325 -4120
rect -1290 -4150 -1220 -4120
rect -1185 -4150 -1125 -4120
rect -2230 -4160 -1125 -4150
rect -2230 -4175 -2180 -4160
rect -2125 -4175 -2075 -4160
rect -2020 -4175 -1970 -4160
rect -1915 -4175 -1865 -4160
rect -1810 -4175 -1760 -4160
rect -1595 -4175 -1545 -4160
rect -1490 -4175 -1440 -4160
rect -1385 -4175 -1335 -4160
rect -1280 -4175 -1230 -4160
rect -1175 -4175 -1125 -4160
rect -1070 -4175 -1020 -4085
rect -2335 -5390 -2285 -5375
rect -2230 -5390 -2180 -5375
rect -2125 -5390 -2075 -5375
rect -2020 -5390 -1970 -5375
rect -1915 -5390 -1865 -5375
rect -1810 -5390 -1760 -5375
rect -1595 -5390 -1545 -5375
rect -1490 -5390 -1440 -5375
rect -1385 -5390 -1335 -5375
rect -1280 -5390 -1230 -5375
rect -1175 -5390 -1125 -5375
rect -1070 -5390 -1020 -5375
<< polycont >>
rect -2165 -145 -2130 -115
rect -2060 -145 -2025 -115
rect -1955 -145 -1920 -115
rect -1745 -145 -1710 -115
rect -1425 -145 -1390 -115
rect -1320 -145 -1285 -115
rect -1215 -145 -1180 -115
rect -2370 -200 -2340 -170
rect -1115 -220 -1085 -190
rect -2430 -1675 -2400 -1645
rect -1145 -2150 -1115 -2120
rect -2325 -2720 -2295 -2690
rect -2375 -4095 -2345 -4065
rect -1120 -4075 -1090 -4045
rect -2170 -4150 -2135 -4120
rect -2065 -4150 -2030 -4120
rect -1960 -4150 -1925 -4120
rect -1750 -4150 -1715 -4120
rect -1430 -4150 -1395 -4120
rect -1325 -4150 -1290 -4120
rect -1220 -4150 -1185 -4120
<< locali >>
rect -2470 1230 -965 1275
rect -2470 1205 -2335 1230
rect -2380 1095 -2335 1205
rect -2380 -75 -2370 1095
rect -2345 -75 -2335 1095
rect -2380 -160 -2335 -75
rect -2275 1150 -1070 1195
rect -2275 1095 -2230 1150
rect -2275 -75 -2265 1095
rect -2240 -75 -2230 1095
rect -2275 -85 -2230 -75
rect -2170 1095 -2125 1105
rect -2170 -75 -2160 1095
rect -2135 -75 -2125 1095
rect -2170 -105 -2125 -75
rect -2065 1095 -2020 1105
rect -2065 -75 -2055 1095
rect -2030 -75 -2020 1095
rect -2065 -105 -2020 -75
rect -1960 1095 -1915 1105
rect -1960 -75 -1950 1095
rect -1925 -75 -1915 1095
rect -1960 -105 -1915 -75
rect -1855 1095 -1810 1150
rect -1855 -75 -1845 1095
rect -1820 -75 -1810 1095
rect -1855 -85 -1810 -75
rect -1750 1095 -1595 1105
rect -1750 -75 -1740 1095
rect -1715 -75 -1685 1095
rect -1660 -75 -1630 1095
rect -1605 -75 -1595 1095
rect -1750 -85 -1595 -75
rect -1535 1095 -1490 1150
rect -1535 -75 -1525 1095
rect -1500 -75 -1490 1095
rect -1535 -85 -1490 -75
rect -1430 1095 -1385 1105
rect -1430 -75 -1420 1095
rect -1395 -75 -1385 1095
rect -1430 -105 -1385 -75
rect -1325 1095 -1280 1105
rect -1325 -75 -1315 1095
rect -1290 -75 -1280 1095
rect -1325 -105 -1280 -75
rect -1220 1095 -1175 1105
rect -1220 -75 -1210 1095
rect -1185 -75 -1175 1095
rect -1220 -105 -1175 -75
rect -1115 1095 -1070 1150
rect -1115 -75 -1105 1095
rect -1080 -75 -1070 1095
rect -1115 -85 -1070 -75
rect -1010 1095 -965 1230
rect -1010 -75 -1000 1095
rect -975 -75 -965 1095
rect -2175 -115 -2120 -105
rect -2175 -145 -2165 -115
rect -2130 -145 -2120 -115
rect -2175 -155 -2120 -145
rect -2070 -115 -2015 -105
rect -2070 -145 -2060 -115
rect -2025 -145 -2015 -115
rect -2070 -155 -2015 -145
rect -1965 -115 -1910 -105
rect -1965 -145 -1955 -115
rect -1920 -145 -1910 -115
rect -1965 -155 -1910 -145
rect -1755 -115 -1700 -105
rect -1755 -145 -1745 -115
rect -1710 -145 -1700 -115
rect -1755 -155 -1700 -145
rect -1435 -115 -1380 -105
rect -1435 -145 -1425 -115
rect -1390 -145 -1380 -115
rect -1435 -155 -1380 -145
rect -1330 -115 -1275 -105
rect -1330 -145 -1320 -115
rect -1285 -145 -1275 -115
rect -1330 -155 -1275 -145
rect -1225 -115 -1170 -105
rect -1225 -145 -1215 -115
rect -1180 -145 -1170 -115
rect -1225 -155 -1170 -145
rect -2380 -170 -2330 -160
rect -2380 -200 -2370 -170
rect -2340 -200 -2330 -170
rect -1755 -175 -1710 -155
rect -2380 -210 -2330 -200
rect -2380 -285 -2335 -210
rect -1870 -220 -1710 -175
rect -1125 -185 -1075 -180
rect -1010 -185 -965 -75
rect -1250 -190 -965 -185
rect -1250 -220 -1115 -190
rect -1085 -220 -965 -190
rect -2380 -1455 -2370 -285
rect -2345 -1455 -2335 -285
rect -2380 -1465 -2335 -1455
rect -2275 -285 -2230 -275
rect -2275 -1455 -2265 -285
rect -2240 -1455 -2230 -285
rect -2275 -1465 -2230 -1455
rect -1870 -285 -1825 -220
rect -1250 -230 -965 -220
rect -1870 -1455 -1860 -285
rect -1835 -1455 -1825 -285
rect -1870 -1465 -1825 -1455
rect -1465 -285 -1310 -275
rect -1465 -1455 -1455 -285
rect -1430 -1455 -1400 -285
rect -1375 -1455 -1345 -285
rect -1320 -1455 -1310 -285
rect -1465 -1465 -1310 -1455
rect -1250 -285 -1205 -230
rect -1250 -1455 -1240 -285
rect -1215 -1455 -1205 -285
rect -1250 -1465 -1205 -1455
rect -2470 -1635 -2425 -1525
rect -2470 -1645 -1175 -1635
rect -2470 -1675 -2430 -1645
rect -2400 -1670 -2355 -1645
rect -1185 -1670 -1175 -1645
rect -2400 -1675 -1175 -1670
rect -2470 -1680 -1175 -1675
rect -2470 -1685 -2390 -1680
rect -2365 -1750 -1175 -1740
rect -2365 -1775 -2355 -1750
rect -1185 -1775 -1175 -1750
rect -2365 -1805 -1175 -1775
rect -2365 -1830 -2355 -1805
rect -1185 -1830 -1175 -1805
rect -2365 -1860 -1175 -1830
rect -2365 -1885 -2355 -1860
rect -1185 -1885 -1175 -1860
rect -2365 -1895 -1175 -1885
rect -2470 -1965 -1175 -1955
rect -2470 -1990 -2355 -1965
rect -1185 -1990 -1175 -1965
rect -2470 -2000 -1175 -1990
rect -2470 -2275 -2425 -2000
rect -2365 -2070 -1175 -2060
rect -2365 -2095 -2355 -2070
rect -1185 -2095 -1175 -2070
rect -2365 -2105 -1175 -2095
rect -1155 -2120 -1105 -2110
rect -1155 -2150 -1145 -2120
rect -1115 -2150 -1105 -2120
rect -1155 -2165 -1105 -2150
rect -2365 -2175 -1105 -2165
rect -2365 -2200 -2355 -2175
rect -1185 -2200 -1105 -2175
rect -2365 -2210 -1105 -2200
rect -2470 -2285 -1175 -2275
rect -2470 -2310 -2355 -2285
rect -1185 -2310 -1175 -2285
rect -2470 -2320 -1175 -2310
rect -2470 -2595 -2425 -2320
rect -2365 -2390 -1175 -2380
rect -2365 -2415 -2355 -2390
rect -1185 -2415 -1175 -2390
rect -2365 -2445 -1175 -2415
rect -2365 -2470 -2355 -2445
rect -1185 -2470 -1175 -2445
rect -2365 -2500 -1175 -2470
rect -2365 -2525 -2355 -2500
rect -1185 -2525 -1175 -2500
rect -2365 -2535 -1175 -2525
rect -2470 -2605 -1175 -2595
rect -2470 -2630 -2355 -2605
rect -1185 -2630 -1175 -2605
rect -2470 -2640 -1175 -2630
rect -2470 -2680 -2425 -2640
rect -2470 -2690 -2285 -2680
rect -2470 -2720 -2325 -2690
rect -2295 -2720 -2285 -2690
rect -2470 -2725 -2285 -2720
rect -2335 -2730 -2285 -2725
rect -2385 -2810 -2340 -2800
rect -2385 -3980 -2375 -2810
rect -2350 -3980 -2340 -2810
rect -2385 -4055 -2340 -3980
rect -2280 -2810 -2235 -2800
rect -2280 -3980 -2270 -2810
rect -2245 -3980 -2235 -2810
rect -2280 -3990 -2235 -3980
rect -1875 -2810 -1830 -2800
rect -1875 -3980 -1865 -2810
rect -1840 -3980 -1830 -2810
rect -1875 -4045 -1830 -3980
rect -1470 -2810 -1315 -2800
rect -1470 -3980 -1460 -2810
rect -1435 -3980 -1405 -2810
rect -1380 -3980 -1350 -2810
rect -1325 -3980 -1315 -2810
rect -1470 -3990 -1315 -3980
rect -1255 -2810 -1210 -2800
rect -1255 -3980 -1245 -2810
rect -1220 -3980 -1210 -2810
rect -1255 -4035 -1210 -3980
rect -1255 -4045 -970 -4035
rect -2385 -4065 -2335 -4055
rect -2385 -4095 -2375 -4065
rect -2345 -4095 -2335 -4065
rect -1875 -4090 -1715 -4045
rect -1255 -4075 -1120 -4045
rect -1090 -4075 -970 -4045
rect -1255 -4080 -970 -4075
rect -1130 -4085 -1080 -4080
rect -2385 -4105 -2335 -4095
rect -2385 -4190 -2340 -4105
rect -1760 -4110 -1715 -4090
rect -2180 -4120 -2125 -4110
rect -2180 -4150 -2170 -4120
rect -2135 -4150 -2125 -4120
rect -2180 -4160 -2125 -4150
rect -2075 -4120 -2020 -4110
rect -2075 -4150 -2065 -4120
rect -2030 -4150 -2020 -4120
rect -2075 -4160 -2020 -4150
rect -1970 -4120 -1915 -4110
rect -1970 -4150 -1960 -4120
rect -1925 -4150 -1915 -4120
rect -1970 -4160 -1915 -4150
rect -1760 -4120 -1705 -4110
rect -1760 -4150 -1750 -4120
rect -1715 -4150 -1705 -4120
rect -1760 -4160 -1705 -4150
rect -1440 -4120 -1385 -4110
rect -1440 -4150 -1430 -4120
rect -1395 -4150 -1385 -4120
rect -1440 -4160 -1385 -4150
rect -1335 -4120 -1280 -4110
rect -1335 -4150 -1325 -4120
rect -1290 -4150 -1280 -4120
rect -1335 -4160 -1280 -4150
rect -1230 -4120 -1175 -4110
rect -1230 -4150 -1220 -4120
rect -1185 -4150 -1175 -4120
rect -1230 -4160 -1175 -4150
rect -2385 -5360 -2375 -4190
rect -2350 -5360 -2340 -4190
rect -2385 -5465 -2340 -5360
rect -2280 -4190 -2235 -4180
rect -2280 -5360 -2270 -4190
rect -2245 -5360 -2235 -4190
rect -2280 -5415 -2235 -5360
rect -2175 -4190 -2130 -4160
rect -2175 -5360 -2165 -4190
rect -2140 -5360 -2130 -4190
rect -2175 -5370 -2130 -5360
rect -2070 -4190 -2025 -4160
rect -2070 -5360 -2060 -4190
rect -2035 -5360 -2025 -4190
rect -2070 -5370 -2025 -5360
rect -1965 -4190 -1920 -4160
rect -1965 -5360 -1955 -4190
rect -1930 -5360 -1920 -4190
rect -1965 -5370 -1920 -5360
rect -1860 -4190 -1815 -4180
rect -1860 -5360 -1850 -4190
rect -1825 -5360 -1815 -4190
rect -1860 -5415 -1815 -5360
rect -1755 -4190 -1600 -4180
rect -1755 -5360 -1745 -4190
rect -1720 -5360 -1690 -4190
rect -1665 -5360 -1635 -4190
rect -1610 -5360 -1600 -4190
rect -1755 -5370 -1600 -5360
rect -1540 -4190 -1495 -4180
rect -1540 -5360 -1530 -4190
rect -1505 -5360 -1495 -4190
rect -1540 -5415 -1495 -5360
rect -1435 -4190 -1390 -4160
rect -1435 -5360 -1425 -4190
rect -1400 -5360 -1390 -4190
rect -1435 -5370 -1390 -5360
rect -1330 -4190 -1285 -4160
rect -1330 -5360 -1320 -4190
rect -1295 -5360 -1285 -4190
rect -1330 -5370 -1285 -5360
rect -1225 -4190 -1180 -4160
rect -1225 -5360 -1215 -4190
rect -1190 -5360 -1180 -4190
rect -1225 -5370 -1180 -5360
rect -1120 -4190 -1075 -4180
rect -1120 -5360 -1110 -4190
rect -1085 -5360 -1075 -4190
rect -1120 -5415 -1075 -5360
rect -2280 -5460 -1075 -5415
rect -1015 -4190 -970 -4080
rect -1015 -5360 -1005 -4190
rect -980 -5360 -970 -4190
rect -2470 -5495 -2340 -5465
rect -1015 -5495 -970 -5360
rect -2470 -5540 -970 -5495
<< viali >>
rect -1740 300 -1715 905
rect -1685 300 -1660 905
rect -1630 300 -1605 905
rect -2265 -1125 -2240 -440
rect -1455 -1125 -1430 -440
rect -1400 -1125 -1375 -440
rect -1345 -1125 -1320 -440
rect -2355 -1775 -1185 -1750
rect -2355 -1830 -1185 -1805
rect -2355 -1885 -1185 -1860
rect -2355 -2095 -1185 -2070
rect -2355 -2415 -1185 -2390
rect -2355 -2470 -1185 -2445
rect -2355 -2525 -1185 -2500
rect -2270 -3730 -2245 -3040
rect -1460 -3730 -1435 -3040
rect -1405 -3730 -1380 -3040
rect -1350 -3730 -1325 -3040
rect -1745 -5090 -1720 -4475
rect -1690 -5090 -1665 -4475
rect -1635 -5090 -1610 -4475
<< metal1 >>
rect -2470 905 -910 920
rect -2470 300 -1740 905
rect -1715 300 -1685 905
rect -1660 300 -1630 905
rect -1605 300 -910 905
rect -2470 295 -910 300
rect -2470 -440 -910 -430
rect -2470 -1125 -2265 -440
rect -2240 -1125 -1455 -440
rect -1430 -1125 -1400 -440
rect -1375 -1125 -1345 -440
rect -1320 -1125 -910 -440
rect -2470 -1130 -910 -1125
rect -2470 -1750 -910 -1735
rect -2470 -1775 -2355 -1750
rect -1185 -1775 -910 -1750
rect -2470 -1805 -910 -1775
rect -2470 -1830 -2355 -1805
rect -1185 -1830 -910 -1805
rect -2470 -1860 -910 -1830
rect -2470 -1885 -2355 -1860
rect -1185 -1885 -910 -1860
rect -2470 -2070 -910 -1885
rect -2470 -2095 -2355 -2070
rect -1185 -2095 -910 -2070
rect -2470 -2160 -910 -2095
rect -2470 -2390 -910 -2375
rect -2470 -2415 -2355 -2390
rect -1185 -2415 -910 -2390
rect -2470 -2445 -910 -2415
rect -2470 -2470 -2355 -2445
rect -1185 -2470 -910 -2445
rect -2470 -2500 -910 -2470
rect -2470 -2525 -2355 -2500
rect -1185 -2525 -910 -2500
rect -2470 -2540 -910 -2525
rect -2470 -3040 -910 -3035
rect -2470 -3730 -2270 -3040
rect -2245 -3730 -1460 -3040
rect -1435 -3730 -1405 -3040
rect -1380 -3730 -1350 -3040
rect -1325 -3730 -910 -3040
rect -2470 -3735 -910 -3730
rect -2470 -4475 -910 -4470
rect -2470 -5090 -1745 -4475
rect -1720 -5090 -1690 -4475
rect -1665 -5090 -1635 -4475
rect -1610 -5090 -910 -4475
rect -2470 -5095 -910 -5090
<< labels >>
rlabel metal1 -2470 -4810 -2470 -4810 7 GND
rlabel metal1 -2470 -3405 -2470 -3405 7 VDD
rlabel locali -2470 -2705 -2470 -2705 7 VBP
rlabel metal1 -2470 -2465 -2470 -2465 7 VDD
rlabel metal1 -2470 -1825 -2470 -1825 7 GND
rlabel locali -2470 -1615 -2470 -1615 7 VBN
rlabel metal1 -2470 -780 -2470 -780 7 GND
rlabel metal1 -2470 530 -2470 530 7 VDD
rlabel locali -2470 1240 -2470 1240 7 VCP
rlabel locali -2470 -5505 -2470 -5505 7 VCN
<< end >>
