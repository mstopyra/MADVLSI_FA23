magic
tech sky130A
timestamp 1694477420
<< nwell >>
rect -125 140 80 280
<< nmos >>
rect -5 -5 10 95
<< pmos >>
rect -5 160 10 260
<< ndiff >>
rect -55 80 -5 95
rect -55 10 -40 80
rect -20 10 -5 80
rect -55 -5 -5 10
rect 10 80 60 95
rect 10 10 25 80
rect 45 10 60 80
rect 10 -5 60 10
<< pdiff >>
rect -55 245 -5 260
rect -55 175 -40 245
rect -20 175 -5 245
rect -55 160 -5 175
rect 10 245 60 260
rect 10 175 25 245
rect 45 175 60 245
rect 10 160 60 175
<< ndiffc >>
rect -40 10 -20 80
rect 25 10 45 80
<< pdiffc >>
rect -40 175 -20 245
rect 25 175 45 245
<< psubdiff >>
rect -105 80 -55 95
rect -105 10 -90 80
rect -70 10 -55 80
rect -105 -5 -55 10
<< nsubdiff >>
rect -105 245 -55 260
rect -105 175 -90 245
rect -70 175 -55 245
rect -105 160 -55 175
<< psubdiffcont >>
rect -90 10 -70 80
<< nsubdiffcont >>
rect -90 175 -70 245
<< poly >>
rect -5 260 10 275
rect -5 95 10 160
rect -5 -20 10 -5
rect -30 -30 10 -20
rect -30 -50 -20 -30
rect 0 -50 10 -30
rect -30 -60 10 -50
<< polycont >>
rect -20 -50 0 -30
<< locali >>
rect -100 245 -10 255
rect -100 175 -90 245
rect -70 175 -40 245
rect -20 175 -10 245
rect -100 165 -10 175
rect 15 245 55 255
rect 15 175 25 245
rect 45 175 55 245
rect 15 165 55 175
rect 35 90 55 165
rect -100 80 -10 90
rect -100 10 -90 80
rect -70 10 -40 80
rect -20 10 -10 80
rect -100 0 -10 10
rect 15 80 55 90
rect 15 10 25 80
rect 45 10 55 80
rect 15 0 55 10
rect 35 -20 55 0
rect -125 -30 10 -20
rect -125 -40 -20 -30
rect -30 -50 -20 -40
rect 0 -50 10 -30
rect 35 -40 80 -20
rect -30 -60 10 -50
<< viali >>
rect -90 175 -70 245
rect -40 175 -20 245
rect -90 10 -70 80
rect -40 10 -20 80
<< metal1 >>
rect -125 245 80 255
rect -125 175 -90 245
rect -70 175 -40 245
rect -20 175 80 245
rect -125 165 80 175
rect -125 80 80 90
rect -125 10 -90 80
rect -70 10 -40 80
rect -20 10 80 80
rect -125 0 80 10
<< labels >>
rlabel metal1 -125 210 -125 210 7 VP
port 3 w
rlabel locali -125 -30 -125 -30 7 A
port 1 w
rlabel locali 80 -30 80 -30 3 Y
port 2 e
rlabel metal1 -125 45 -125 45 7 VN
port 4 w
<< end >>
