magic
tech sky130A
timestamp 1695926555
<< nwell >>
rect -445 335 155 805
<< nmos >>
rect -375 -115 -360 285
rect -145 170 -130 270
rect -80 170 -65 270
rect -15 170 0 270
rect -145 -35 -130 65
rect -80 -35 -65 65
rect -15 -35 0 65
<< pmos >>
rect -375 630 -360 730
rect -310 630 -295 730
rect -375 355 -360 455
rect -310 355 -295 455
rect -120 385 -105 785
rect 5 630 20 730
rect 25 420 40 520
<< ndiff >>
rect -425 80 -375 285
rect -425 -90 -410 80
rect -390 -90 -375 80
rect -425 -115 -375 -90
rect -360 80 -310 285
rect -195 255 -145 270
rect -195 185 -180 255
rect -160 185 -145 255
rect -195 170 -145 185
rect -130 255 -80 270
rect -130 185 -115 255
rect -95 185 -80 255
rect -130 170 -80 185
rect -65 255 -15 270
rect -65 185 -50 255
rect -30 185 -15 255
rect -65 170 -15 185
rect 0 255 50 270
rect 0 185 15 255
rect 35 185 50 255
rect 0 170 50 185
rect -360 -90 -345 80
rect -325 -90 -310 80
rect -195 50 -145 65
rect -195 -20 -180 50
rect -160 -20 -145 50
rect -195 -35 -145 -20
rect -130 50 -80 65
rect -130 -20 -115 50
rect -95 -20 -80 50
rect -130 -35 -80 -20
rect -65 50 -15 65
rect -65 -20 -50 50
rect -30 -20 -15 50
rect -65 -35 -15 -20
rect 0 50 50 65
rect 0 -20 15 50
rect 35 -20 50 50
rect 0 -35 50 -20
rect -360 -115 -310 -90
<< pdiff >>
rect -170 770 -120 785
rect -425 715 -375 730
rect -425 645 -410 715
rect -390 645 -375 715
rect -425 630 -375 645
rect -360 715 -310 730
rect -360 645 -345 715
rect -325 645 -310 715
rect -360 630 -310 645
rect -295 715 -245 730
rect -295 645 -280 715
rect -260 645 -245 715
rect -295 630 -245 645
rect -170 600 -155 770
rect -135 600 -120 770
rect -425 440 -375 455
rect -425 370 -410 440
rect -390 370 -375 440
rect -425 355 -375 370
rect -360 440 -310 455
rect -360 370 -345 440
rect -325 370 -310 440
rect -360 355 -310 370
rect -295 440 -245 455
rect -295 370 -280 440
rect -260 370 -245 440
rect -170 385 -120 600
rect -105 770 -55 785
rect -105 600 -90 770
rect -70 730 -55 770
rect -70 715 5 730
rect -70 645 -30 715
rect -10 645 5 715
rect -70 630 5 645
rect 20 715 70 730
rect 20 645 35 715
rect 55 645 70 715
rect 20 630 70 645
rect -70 600 -55 630
rect -105 385 -55 600
rect -25 505 25 520
rect -25 435 -10 505
rect 10 435 25 505
rect -25 420 25 435
rect 40 505 90 520
rect 40 435 55 505
rect 75 435 90 505
rect 40 420 90 435
rect -295 355 -245 370
<< ndiffc >>
rect -410 -90 -390 80
rect -180 185 -160 255
rect -115 185 -95 255
rect -50 185 -30 255
rect 15 185 35 255
rect -345 -90 -325 80
rect -180 -20 -160 50
rect -115 -20 -95 50
rect -50 -20 -30 50
rect 15 -20 35 50
<< pdiffc >>
rect -410 645 -390 715
rect -345 645 -325 715
rect -280 645 -260 715
rect -155 600 -135 770
rect -410 370 -390 440
rect -345 370 -325 440
rect -280 370 -260 440
rect -90 600 -70 770
rect -30 645 -10 715
rect 35 645 55 715
rect -10 435 10 505
rect 55 435 75 505
<< psubdiff >>
rect 50 50 100 65
rect 50 -20 65 50
rect 85 -20 100 50
rect 50 -35 100 -20
<< nsubdiff >>
rect -245 715 -200 730
rect -245 645 -235 715
rect -215 645 -200 715
rect -245 630 -200 645
<< psubdiffcont >>
rect 65 -20 85 50
<< nsubdiffcont >>
rect -235 645 -215 715
<< poly >>
rect -120 785 -105 800
rect -375 730 -360 745
rect -310 730 -295 745
rect -375 455 -360 630
rect -310 615 -295 630
rect -310 605 -230 615
rect -310 600 -265 605
rect -275 580 -265 600
rect -240 580 -230 605
rect -275 570 -230 580
rect -335 545 -290 555
rect -335 520 -325 545
rect -300 520 -290 545
rect -335 510 -290 520
rect -335 480 -320 510
rect -335 465 -295 480
rect -310 455 -295 465
rect 5 730 20 745
rect 5 610 20 630
rect -40 600 20 610
rect -40 575 -30 600
rect -5 595 20 600
rect 95 595 140 605
rect -5 575 5 595
rect -40 565 5 575
rect 95 570 105 595
rect 130 570 140 595
rect 95 560 140 570
rect 95 545 110 560
rect 25 530 110 545
rect 25 520 40 530
rect 25 405 40 420
rect -20 395 40 405
rect -120 375 -105 385
rect -215 360 -170 370
rect -120 360 -65 375
rect -20 370 -10 395
rect 15 390 40 395
rect 15 370 25 390
rect -20 360 25 370
rect -375 285 -360 355
rect -310 340 -295 355
rect -215 340 -205 360
rect -310 335 -205 340
rect -180 335 -170 360
rect -310 325 -170 335
rect -295 290 -130 300
rect -295 265 -285 290
rect -260 285 -130 290
rect -260 265 -250 285
rect -295 255 -250 265
rect -225 165 -210 285
rect -145 270 -130 285
rect -80 270 -65 360
rect 30 320 75 330
rect 30 300 40 320
rect -15 295 40 300
rect 65 300 75 320
rect 65 295 125 300
rect -15 285 125 295
rect -15 270 0 285
rect -255 155 -210 165
rect -145 155 -130 170
rect -255 130 -245 155
rect -220 130 -210 155
rect -255 120 -210 130
rect -150 115 -105 125
rect -150 90 -140 115
rect -115 90 -105 115
rect -150 80 -105 90
rect -145 65 -130 80
rect -80 65 -65 170
rect -15 155 0 170
rect -40 115 5 125
rect -40 90 -30 115
rect -5 90 5 115
rect -40 80 5 90
rect -15 65 0 80
rect -145 -50 -130 -35
rect -445 -135 -400 -125
rect -375 -135 -360 -115
rect -80 -135 -65 -35
rect -15 -50 0 -35
rect 110 -75 125 285
rect -40 -85 125 -75
rect -40 -110 -30 -85
rect -5 -90 125 -85
rect -5 -110 5 -90
rect -40 -120 5 -110
rect -445 -160 -435 -135
rect -410 -150 -65 -135
rect -410 -160 -400 -150
rect -445 -170 -400 -160
<< polycont >>
rect -265 580 -240 605
rect -325 520 -300 545
rect -30 575 -5 600
rect 105 570 130 595
rect -10 370 15 395
rect -205 335 -180 360
rect -285 265 -260 290
rect 40 295 65 320
rect -245 130 -220 155
rect -140 90 -115 115
rect -30 90 -5 115
rect -30 -110 -5 -85
rect -435 -160 -410 -135
<< locali >>
rect -165 770 -125 780
rect -165 725 -155 770
rect -420 715 -380 725
rect -420 645 -410 715
rect -390 645 -380 715
rect -420 605 -380 645
rect -445 560 -380 605
rect -355 715 -315 725
rect -355 645 -345 715
rect -325 645 -315 715
rect -355 635 -315 645
rect -290 715 -155 725
rect -290 645 -280 715
rect -260 645 -235 715
rect -215 645 -155 715
rect -290 635 -155 645
rect -355 575 -335 635
rect -275 605 -230 615
rect -275 580 -265 605
rect -240 580 -230 605
rect -165 600 -155 635
rect -135 600 -125 770
rect -165 590 -125 600
rect -100 770 -60 780
rect -100 600 -90 770
rect -70 725 -60 770
rect -70 715 0 725
rect -70 645 -30 715
rect -10 645 0 715
rect -70 635 0 645
rect 25 715 65 725
rect 25 645 35 715
rect 55 645 65 715
rect 25 635 65 645
rect -70 600 -60 635
rect -100 590 -60 600
rect -40 600 5 610
rect -355 555 -315 575
rect -275 570 -230 580
rect -335 545 -290 555
rect -335 520 -325 545
rect -300 520 -290 545
rect -335 510 -290 520
rect -265 490 -245 570
rect -335 470 -245 490
rect -335 450 -315 470
rect -155 450 -135 590
rect -90 515 -70 590
rect -40 575 -30 600
rect -5 575 5 600
rect 45 605 65 635
rect 45 595 155 605
rect 45 585 105 595
rect -40 565 5 575
rect 95 570 105 585
rect 130 570 155 595
rect -15 545 70 565
rect 95 560 155 570
rect 45 515 70 545
rect -90 505 20 515
rect -90 495 -10 505
rect -420 440 -380 450
rect -420 405 -410 440
rect -445 370 -410 405
rect -390 370 -380 440
rect -445 360 -380 370
rect -355 440 -315 450
rect -355 370 -345 440
rect -325 370 -315 440
rect -355 360 -315 370
rect -290 440 -135 450
rect -290 370 -280 440
rect -260 430 -135 440
rect -20 435 -10 495
rect 10 435 20 505
rect -260 370 -250 430
rect -20 425 20 435
rect 45 505 85 515
rect 45 435 55 505
rect 75 435 85 505
rect 45 425 85 435
rect 55 405 75 425
rect -20 395 25 405
rect -20 380 -10 395
rect -40 370 -10 380
rect 15 370 25 395
rect -290 360 -250 370
rect -215 360 -170 370
rect -335 275 -315 360
rect -215 335 -205 360
rect -180 345 -170 360
rect -40 360 25 370
rect 55 360 155 405
rect -180 335 -105 345
rect -215 325 -105 335
rect -295 290 -250 300
rect -295 275 -285 290
rect -335 265 -285 275
rect -260 265 -250 290
rect -125 265 -105 325
rect -40 265 -20 360
rect 55 330 75 360
rect 30 320 75 330
rect 30 295 40 320
rect 65 295 75 320
rect 30 285 75 295
rect -335 255 -250 265
rect -190 255 -150 265
rect -190 225 -180 255
rect -295 205 -180 225
rect -295 90 -275 205
rect -190 185 -180 205
rect -160 185 -150 255
rect -190 175 -150 185
rect -125 255 -85 265
rect -125 185 -115 255
rect -95 185 -85 255
rect -125 175 -85 185
rect -60 255 -20 265
rect -60 185 -50 255
rect -30 185 -20 255
rect -60 175 -20 185
rect 5 255 45 265
rect 5 185 15 255
rect 35 185 45 255
rect 5 175 45 185
rect -255 155 -210 165
rect -255 130 -245 155
rect -220 130 -210 155
rect -255 120 -210 130
rect -420 80 -380 90
rect -420 -90 -410 80
rect -390 -90 -380 80
rect -420 -100 -380 -90
rect -355 80 -275 90
rect -355 -90 -345 80
rect -325 70 -275 80
rect -325 -90 -315 70
rect -230 -55 -210 120
rect -190 60 -170 175
rect -125 125 -105 175
rect -150 115 -105 125
rect -150 90 -140 115
rect -115 90 -105 115
rect -150 80 -105 90
rect -40 125 -20 175
rect -40 115 5 125
rect -40 90 -30 115
rect -5 90 5 115
rect 25 110 45 175
rect 25 90 95 110
rect -40 80 5 90
rect 75 60 95 90
rect -190 50 -150 60
rect -190 -20 -180 50
rect -160 -20 -150 50
rect -190 -30 -150 -20
rect -125 50 -85 60
rect -125 -20 -115 50
rect -95 -20 -85 50
rect -125 -30 -85 -20
rect -60 50 -20 60
rect -60 -20 -50 50
rect -30 -20 -20 50
rect -60 -30 -20 -20
rect 5 50 95 60
rect 5 -20 15 50
rect 35 -20 65 50
rect 85 -20 95 50
rect 5 -30 95 -20
rect -125 -55 -105 -30
rect -230 -75 -105 -55
rect -40 -75 -20 -30
rect -355 -100 -315 -90
rect -40 -85 5 -75
rect -40 -110 -30 -85
rect -5 -110 5 -85
rect -40 -120 5 -110
rect -445 -135 -400 -125
rect -445 -160 -435 -135
rect -410 -160 -400 -135
rect -445 -170 -400 -160
<< viali >>
rect -280 645 -260 715
rect -235 645 -215 715
rect -410 -90 -390 80
rect 15 -20 35 50
rect 65 -20 85 50
rect -435 -160 -410 -135
<< metal1 >>
rect -445 715 155 725
rect -445 645 -280 715
rect -260 645 -235 715
rect -215 645 155 715
rect -445 635 155 645
rect -445 80 155 90
rect -445 -90 -410 80
rect -390 50 155 80
rect -390 -20 15 50
rect 35 -20 65 50
rect 85 -20 155 50
rect -390 -90 155 -20
rect -445 -100 155 -90
rect -445 -135 155 -125
rect -445 -160 -435 -135
rect -410 -160 155 -135
rect -445 -170 155 -160
<< labels >>
rlabel metal1 -445 680 -445 680 7 VDD
rlabel locali -445 580 -445 580 7 D
rlabel locali -445 380 -445 380 7 DB
rlabel metal1 -445 -10 -445 -10 7 GND
rlabel metal1 -445 -150 -445 -150 7 CLK
rlabel locali 155 580 155 580 3 Q
rlabel locali 155 380 155 380 3 QB
<< end >>
