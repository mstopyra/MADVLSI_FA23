magic
tech sky130A
timestamp 1697753258
<< nwell >>
rect -840 7060 -460 7110
rect -345 7065 1410 7110
rect -510 6855 -460 7060
rect -395 6855 1410 7065
rect -510 6805 1410 6855
rect -395 5830 1410 6805
rect -345 5640 1410 5830
<< poly >>
rect -840 7060 -460 7110
rect -510 6855 -460 7060
rect -510 6845 -215 6855
rect -510 6815 -255 6845
rect -225 6815 -215 6845
rect -510 6805 -215 6815
rect -265 5605 -215 5615
rect -265 5575 -255 5605
rect -225 5575 -215 5605
rect -265 5390 -215 5575
rect -265 5360 -255 5390
rect -225 5360 -215 5390
rect -265 5350 -215 5360
<< polycont >>
rect -255 6815 -225 6845
rect -255 5575 -225 5605
rect -255 5360 -225 5390
<< locali >>
rect -395 6995 -150 7065
rect -395 5830 -345 6995
rect -265 6845 -215 6855
rect -265 6815 -255 6845
rect -225 6815 -215 6845
rect -265 5605 -215 6815
rect -265 5575 -255 5605
rect -225 5575 -215 5605
rect -265 5565 -215 5575
rect -345 5465 -105 5515
rect -265 5390 -215 5400
rect -265 5360 -255 5390
rect -225 5360 -215 5390
rect -395 325 -345 3900
rect -265 3835 -215 5360
rect -150 4265 -105 5465
rect -265 3780 -130 3835
rect -395 250 -145 325
<< metal1 >>
rect -345 6135 -140 6710
rect 1410 6085 1515 6135
rect -350 4660 -85 5125
rect -540 3675 -115 3710
rect -540 3635 -110 3675
rect -535 3630 -110 3635
rect 1465 3415 1515 6085
rect 1395 3365 1515 3415
rect 1395 3360 1410 3365
rect 1360 3250 1410 3290
rect 1355 2750 1410 3250
use biasgen  biasgen_0
timestamp 1697752574
transform 1 0 2320 0 1 5790
box -2470 -5540 -910 1300
use FCDA  FCDA_0
timestamp 1697751355
transform 1 0 -125 0 1 3345
box -1760 -730 -220 3765
<< end >>
