* NGSPICE file created from biasgen.ext - technology: sky130A


* Top level circuit biasgen

X0 a_n4050_n2940# VBN a_n4200_n2940# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X1 VBP VBN GND GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X2 a_n3090_n2940# VBN a_n3240_n2940# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X3 a_n3900_n2940# VBN a_n4050_n2940# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X4 a_n3240_n2940# VBN a_n3390_n2940# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X5 a_n4460_n10780# a_n4460_n10780# a_n4460_n10780# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=39.6 ps=151 w=12 l=0.5
X6 a_n4450_n310# a_n4450_n310# a_n4450_n310# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=39.6 ps=151 w=12 l=0.5
X7 GND VBN VBN GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=6.6 ps=25.1 w=12 l=0.5
X8 GND VBN VBP GND sky130_fd_pr__nfet_01v8 ad=6.6 pd=25.1 as=3.3 ps=12.6 w=12 l=0.5
X9 a_n4560_n180# VCP VCP VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=6.6 ps=25.1 w=12 l=0.5
X10 VDD VBP VCN VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=6.6 ps=25.1 w=12 l=0.5
X11 a_n3910_n7990# VBP a_n4060_n7990# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X12 VDD VBP a_n3100_n7990# VDD sky130_fd_pr__pfet_01v8 ad=6.6 pd=25.1 as=1.5 ps=12.2 w=12 l=0.5
X13 a_n4460_n10780# VBP a_n3910_n7990# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=1.5 ps=12.2 w=12 l=0.5
X14 a_n4570_n10750# a_n4460_n10780# GND GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=6.6 ps=25.1 w=12 l=0.5
X15 a_n4460_n10780# a_n4460_n10780# a_n4460_n10780# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=0 ps=0 w=12 l=0.5
X16 GND VBN VCP GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=6.6 ps=25.1 w=12 l=0.5
X17 VBN VBN GND GND sky130_fd_pr__nfet_01v8 ad=6.6 pd=25.1 as=6.6 ps=25.1 w=12 l=0.5
X18 a_n4450_n310# a_n4450_n310# a_n4560_n180# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X19 GND VBN a_n3090_n2940# GND sky130_fd_pr__nfet_01v8 ad=6.6 pd=25.1 as=1.5 ps=12.2 w=12 l=0.5
X20 a_n4570_n10750# a_n4460_n10780# a_n4460_n10780# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X21 a_n4450_n310# VBN a_n3900_n2940# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=1.5 ps=12.2 w=12 l=0.5
X22 VCN VBP VDD VDD sky130_fd_pr__pfet_01v8 ad=6.6 pd=25.1 as=6.6 ps=25.1 w=12 l=0.5
X23 VCP VCP a_n4560_n180# VDD sky130_fd_pr__pfet_01v8 ad=6.6 pd=25.1 as=3.3 ps=12.6 w=12 l=0.5
X24 VCN VCN a_n4570_n10750# GND sky130_fd_pr__nfet_01v8 ad=6.6 pd=25.1 as=3.3 ps=12.6 w=12 l=0.5
X25 a_n4450_n310# a_n4450_n310# a_n4450_n310# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=0 ps=0 w=12 l=0.5
X26 a_n4570_n10750# VCN VCN GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=6.6 ps=25.1 w=12 l=0.5
X27 VCP VBN GND GND sky130_fd_pr__nfet_01v8 ad=6.6 pd=25.1 as=6.6 ps=25.1 w=12 l=0.5
X28 a_n4360_n7990# VBP VDD VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=3.3 ps=12.6 w=12 l=0.5
X29 VDD VBP VBP VDD sky130_fd_pr__pfet_01v8 ad=6.6 pd=25.1 as=6.6 ps=25.1 w=12 l=0.5
X30 a_n3400_n7990# VBP a_n3550_n7990# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X31 a_n4570_n10750# a_n4460_n10780# a_n4460_n10780# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X32 a_n4560_n180# a_n4450_n310# a_n4450_n310# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X33 a_n3550_n7990# VBP a_n4460_n10780# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=3.3 ps=12.6 w=12 l=0.5
X34 a_n4460_n10780# a_n4460_n10780# a_n4570_n10750# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X35 a_n4200_n2940# VBN a_n4350_n2940# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X36 a_n4450_n310# a_n4450_n310# a_n4450_n310# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=0 ps=0 w=12 l=0.5
X37 a_n4350_n2940# VBN GND GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=3.3 ps=12.6 w=12 l=0.5
X38 VBP VBP VDD VDD sky130_fd_pr__pfet_01v8 ad=6.6 pd=25.1 as=6.6 ps=25.1 w=12 l=0.5
X39 VDD a_n4450_n310# a_n4560_n180# VDD sky130_fd_pr__pfet_01v8 ad=6.6 pd=25.1 as=3.3 ps=12.6 w=12 l=0.5
X40 GND a_n4460_n10780# a_n4570_n10750# GND sky130_fd_pr__nfet_01v8 ad=6.6 pd=25.1 as=3.3 ps=12.6 w=12 l=0.5
X41 a_n3390_n2940# VBN a_n3540_n2940# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X42 a_n4460_n10780# a_n4460_n10780# a_n4460_n10780# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=0 ps=0 w=12 l=0.5
X43 a_n3540_n2940# VBN a_n4450_n310# GND sky130_fd_pr__nfet_01v8 ad=1.5 pd=12.2 as=3.3 ps=12.6 w=12 l=0.5
X44 a_n4560_n180# a_n4450_n310# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=6.6 ps=25.1 w=12 l=0.5
X45 a_n4060_n7990# VBP a_n4210_n7990# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X46 a_n4450_n310# a_n4450_n310# a_n4450_n310# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=0 ps=0 w=12 l=0.5
X47 a_n4210_n7990# VBP a_n4360_n7990# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X48 a_n3100_n7990# VBP a_n3250_n7990# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X49 a_n4460_n10780# a_n4460_n10780# a_n4460_n10780# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=0 ps=0 w=12 l=0.5
X50 a_n4450_n310# a_n4450_n310# a_n4560_n180# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X51 a_n4560_n180# a_n4450_n310# a_n4450_n310# VDD sky130_fd_pr__pfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
X52 a_n3250_n7990# VBP a_n3400_n7990# VDD sky130_fd_pr__pfet_01v8 ad=1.5 pd=12.2 as=1.5 ps=12.2 w=12 l=0.5
X53 a_n4460_n10780# a_n4460_n10780# a_n4570_n10750# GND sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.6 as=3.3 ps=12.6 w=12 l=0.5
.end

